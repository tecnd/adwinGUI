module DoubleHiThenLo(tenMHz_ext_clk, 