module synclock_divider(int_ref_clock, synclock, SDIO, SCLK);

input 